-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bbb",
     9 => x"dc080b0b",
    10 => x"0bbbe008",
    11 => x"0b0b0bbb",
    12 => x"e4080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"bbe40c0b",
    16 => x"0b0bbbe0",
    17 => x"0c0b0b0b",
    18 => x"bbdc0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb1e8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"bbdc7080",
    57 => x"c68c278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"5188f804",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bbbec0c",
    65 => x"9f0bbbf0",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"bbf008ff",
    69 => x"05bbf00c",
    70 => x"bbf00880",
    71 => x"25eb38bb",
    72 => x"ec08ff05",
    73 => x"bbec0cbb",
    74 => x"ec088025",
    75 => x"d738800b",
    76 => x"bbf00c80",
    77 => x"0bbbec0c",
    78 => x"0284050d",
    79 => x"0402f005",
    80 => x"0df88053",
    81 => x"f8a05483",
    82 => x"bf527370",
    83 => x"81055533",
    84 => x"51707370",
    85 => x"81055534",
    86 => x"ff125271",
    87 => x"8025eb38",
    88 => x"fbc0539f",
    89 => x"52a07370",
    90 => x"81055534",
    91 => x"ff125271",
    92 => x"8025f238",
    93 => x"0290050d",
    94 => x"0402f405",
    95 => x"0d74538e",
    96 => x"0bbbec08",
    97 => x"258f3882",
    98 => x"bd2dbbec",
    99 => x"08ff05bb",
   100 => x"ec0c82ff",
   101 => x"04bbec08",
   102 => x"bbf00853",
   103 => x"51728a2e",
   104 => x"098106b7",
   105 => x"38715171",
   106 => x"9f24a038",
   107 => x"bbec08a0",
   108 => x"2911f880",
   109 => x"115151a0",
   110 => x"7134bbf0",
   111 => x"088105bb",
   112 => x"f00cbbf0",
   113 => x"08519f71",
   114 => x"25e23880",
   115 => x"0bbbf00c",
   116 => x"bbec0881",
   117 => x"05bbec0c",
   118 => x"83ef0470",
   119 => x"a02912f8",
   120 => x"80115151",
   121 => x"727134bb",
   122 => x"f0088105",
   123 => x"bbf00cbb",
   124 => x"f008a02e",
   125 => x"0981068e",
   126 => x"38800bbb",
   127 => x"f00cbbec",
   128 => x"088105bb",
   129 => x"ec0c028c",
   130 => x"050d0402",
   131 => x"e8050d77",
   132 => x"79565688",
   133 => x"0bfc1677",
   134 => x"712c8f06",
   135 => x"54525480",
   136 => x"53727225",
   137 => x"95387153",
   138 => x"fbe01451",
   139 => x"87713481",
   140 => x"14ff1454",
   141 => x"5472f138",
   142 => x"7153f915",
   143 => x"76712c87",
   144 => x"06535171",
   145 => x"802e8b38",
   146 => x"fbe01451",
   147 => x"71713481",
   148 => x"1454728e",
   149 => x"2495388f",
   150 => x"733153fb",
   151 => x"e01451a0",
   152 => x"71348114",
   153 => x"ff145454",
   154 => x"72f13802",
   155 => x"98050d04",
   156 => x"02ec050d",
   157 => x"800bbbf4",
   158 => x"0cf68c08",
   159 => x"f6900871",
   160 => x"882c5654",
   161 => x"81ff0652",
   162 => x"73722588",
   163 => x"38715482",
   164 => x"0bbbf40c",
   165 => x"72882c73",
   166 => x"81ff0654",
   167 => x"55747325",
   168 => x"8b3872bb",
   169 => x"f4088407",
   170 => x"bbf40c55",
   171 => x"73842b86",
   172 => x"a0712583",
   173 => x"7131700b",
   174 => x"0b0bb7a4",
   175 => x"0c81712b",
   176 => x"ff05f688",
   177 => x"0cfdfc13",
   178 => x"ff122c78",
   179 => x"8829ff94",
   180 => x"0570812c",
   181 => x"bbf40852",
   182 => x"58525551",
   183 => x"52547680",
   184 => x"2e853870",
   185 => x"81075170",
   186 => x"f6940c71",
   187 => x"098105f6",
   188 => x"800c7209",
   189 => x"8105f684",
   190 => x"0c029405",
   191 => x"0d0402f4",
   192 => x"050d7453",
   193 => x"72708105",
   194 => x"5480f52d",
   195 => x"5271802e",
   196 => x"89387151",
   197 => x"82f92d86",
   198 => x"8404810b",
   199 => x"bbdc0c02",
   200 => x"8c050d04",
   201 => x"02fc050d",
   202 => x"81808051",
   203 => x"c0115170",
   204 => x"fb380284",
   205 => x"050d0402",
   206 => x"fc050d84",
   207 => x"bf5186a4",
   208 => x"2dff1151",
   209 => x"708025f6",
   210 => x"38028405",
   211 => x"0d0402fc",
   212 => x"050dec51",
   213 => x"83710c86",
   214 => x"a42d8271",
   215 => x"0c028405",
   216 => x"0d0402fc",
   217 => x"050dec51",
   218 => x"80c2710c",
   219 => x"86a42d82",
   220 => x"710c0284",
   221 => x"050d0402",
   222 => x"fc050dec",
   223 => x"5192710c",
   224 => x"86a42d82",
   225 => x"710c0284",
   226 => x"050d0402",
   227 => x"d0050d7d",
   228 => x"54807453",
   229 => x"bbf8525b",
   230 => x"a9872dbb",
   231 => x"dc087b2e",
   232 => x"81af38bb",
   233 => x"fc0870f8",
   234 => x"0c891580",
   235 => x"f52d8a16",
   236 => x"80f52d71",
   237 => x"82802905",
   238 => x"881780f5",
   239 => x"2d708480",
   240 => x"802912f4",
   241 => x"0c575556",
   242 => x"58a40bec",
   243 => x"0c7aff19",
   244 => x"585a767b",
   245 => x"2e8b3881",
   246 => x"1a77812a",
   247 => x"585a76f7",
   248 => x"38f71a5a",
   249 => x"815b8078",
   250 => x"2580e638",
   251 => x"79527651",
   252 => x"848b2dbc",
   253 => x"c452bbf8",
   254 => x"51abc62d",
   255 => x"bbdc0880",
   256 => x"2eb838bc",
   257 => x"c45c83fc",
   258 => x"597b7084",
   259 => x"055d0870",
   260 => x"81ff0671",
   261 => x"882a7081",
   262 => x"ff067390",
   263 => x"2a7081ff",
   264 => x"0675982a",
   265 => x"e80ce80c",
   266 => x"58e80c57",
   267 => x"e80cfc1a",
   268 => x"5a537880",
   269 => x"25d33888",
   270 => x"c104bbdc",
   271 => x"085b8480",
   272 => x"58bbf851",
   273 => x"ab982dfc",
   274 => x"80188118",
   275 => x"585887e6",
   276 => x"0486b72d",
   277 => x"840bec0c",
   278 => x"7a802e8d",
   279 => x"38b7a851",
   280 => x"91ad2d8f",
   281 => x"b02d88ef",
   282 => x"04b9ac51",
   283 => x"91ad2d7a",
   284 => x"bbdc0c02",
   285 => x"b0050d04",
   286 => x"02d4050d",
   287 => x"8055840b",
   288 => x"ec0c8f91",
   289 => x"2d8bfb2d",
   290 => x"81f82d9f",
   291 => x"fc2dbbdc",
   292 => x"08752e82",
   293 => x"d1388c0b",
   294 => x"ec0cb5e4",
   295 => x"52bbf851",
   296 => x"a9872dbb",
   297 => x"dc08752e",
   298 => x"818338bb",
   299 => x"fc0875ff",
   300 => x"12595b58",
   301 => x"76752e8b",
   302 => x"38811a77",
   303 => x"812a585a",
   304 => x"76f738f7",
   305 => x"1a5a8078",
   306 => x"2580e238",
   307 => x"79527651",
   308 => x"848b2dbc",
   309 => x"c452bbf8",
   310 => x"51abc62d",
   311 => x"bbdc0880",
   312 => x"2eb838bc",
   313 => x"c45b83fc",
   314 => x"597a7084",
   315 => x"055c0870",
   316 => x"81ff0671",
   317 => x"882a7081",
   318 => x"ff067390",
   319 => x"2a7081ff",
   320 => x"0675982a",
   321 => x"e80ce80c",
   322 => x"58e80c57",
   323 => x"e80cfc1a",
   324 => x"5a537880",
   325 => x"25d3388a",
   326 => x"9d048480",
   327 => x"58bbf851",
   328 => x"ab982dfc",
   329 => x"80188118",
   330 => x"585889c6",
   331 => x"04bbfc08",
   332 => x"f80c86b7",
   333 => x"2d840bec",
   334 => x"0c878b51",
   335 => x"b1e02db7",
   336 => x"a85191ad",
   337 => x"2d8fb02d",
   338 => x"8c872d91",
   339 => x"bd2db7d4",
   340 => x"0b80f52d",
   341 => x"70822b84",
   342 => x"06b7c80b",
   343 => x"80f52d83",
   344 => x"067107b7",
   345 => x"e00b80f5",
   346 => x"2d70832b",
   347 => x"b806b7ec",
   348 => x"0b80f52d",
   349 => x"70862b80",
   350 => x"c0067473",
   351 => x"0707b7f8",
   352 => x"0b80f52d",
   353 => x"70882b82",
   354 => x"8006b884",
   355 => x"0b80f52d",
   356 => x"70892b84",
   357 => x"80067473",
   358 => x"0707b890",
   359 => x"0b80f52d",
   360 => x"708a2b88",
   361 => x"8006b89c",
   362 => x"0b80f52d",
   363 => x"708c2ba0",
   364 => x"80067473",
   365 => x"0707b8a8",
   366 => x"0b80f52d",
   367 => x"708f2b82",
   368 => x"80800672",
   369 => x"07fc0c53",
   370 => x"54545454",
   371 => x"54545454",
   372 => x"545b5452",
   373 => x"57545486",
   374 => x"53bbdc08",
   375 => x"83388453",
   376 => x"72ec0c8a",
   377 => x"c804800b",
   378 => x"bbdc0c02",
   379 => x"ac050d04",
   380 => x"71980c04",
   381 => x"ffb008bb",
   382 => x"dc0c0481",
   383 => x"0bffb00c",
   384 => x"04800bff",
   385 => x"b00c0402",
   386 => x"f4050d8d",
   387 => x"8904bbdc",
   388 => x"0881f02e",
   389 => x"09810689",
   390 => x"38810bba",
   391 => x"900c8d89",
   392 => x"04bbdc08",
   393 => x"81e02e09",
   394 => x"81068938",
   395 => x"810bba94",
   396 => x"0c8d8904",
   397 => x"bbdc0852",
   398 => x"ba940880",
   399 => x"2e8838bb",
   400 => x"dc088180",
   401 => x"05527184",
   402 => x"2c728f06",
   403 => x"5353ba90",
   404 => x"08802e99",
   405 => x"38728429",
   406 => x"b9d00572",
   407 => x"1381712b",
   408 => x"70097308",
   409 => x"06730c51",
   410 => x"53538cff",
   411 => x"04728429",
   412 => x"b9d00572",
   413 => x"1383712b",
   414 => x"72080772",
   415 => x"0c535380",
   416 => x"0bba940c",
   417 => x"800bba90",
   418 => x"0cbc8451",
   419 => x"8e8a2dbb",
   420 => x"dc08ff24",
   421 => x"fef83880",
   422 => x"0bbbdc0c",
   423 => x"028c050d",
   424 => x"0402f805",
   425 => x"0db9d052",
   426 => x"8f518072",
   427 => x"70840554",
   428 => x"0cff1151",
   429 => x"708025f2",
   430 => x"38028805",
   431 => x"0d0402f0",
   432 => x"050d7551",
   433 => x"8c812d70",
   434 => x"822cfc06",
   435 => x"b9d01172",
   436 => x"109e0671",
   437 => x"0870722a",
   438 => x"70830682",
   439 => x"742b7009",
   440 => x"7406760c",
   441 => x"54515657",
   442 => x"5351538b",
   443 => x"fb2d71bb",
   444 => x"dc0c0290",
   445 => x"050d0402",
   446 => x"fc050d72",
   447 => x"5180710c",
   448 => x"800b8412",
   449 => x"0c028405",
   450 => x"0d0402f0",
   451 => x"050d7570",
   452 => x"08841208",
   453 => x"535353ff",
   454 => x"5471712e",
   455 => x"a8388c81",
   456 => x"2d841308",
   457 => x"70842914",
   458 => x"88117008",
   459 => x"7081ff06",
   460 => x"84180881",
   461 => x"11870684",
   462 => x"1a0c5351",
   463 => x"55515151",
   464 => x"8bfb2d71",
   465 => x"5473bbdc",
   466 => x"0c029005",
   467 => x"0d0402f8",
   468 => x"050d8c81",
   469 => x"2de00870",
   470 => x"8b2a7081",
   471 => x"06515252",
   472 => x"70802e9d",
   473 => x"38bc8408",
   474 => x"708429bc",
   475 => x"8c057381",
   476 => x"ff06710c",
   477 => x"5151bc84",
   478 => x"08811187",
   479 => x"06bc840c",
   480 => x"51800bbc",
   481 => x"ac0c8bf4",
   482 => x"2d8bfb2d",
   483 => x"0288050d",
   484 => x"0402fc05",
   485 => x"0dbc8451",
   486 => x"8df72d8d",
   487 => x"a12d8ece",
   488 => x"518bf02d",
   489 => x"0284050d",
   490 => x"04bcb008",
   491 => x"bbdc0c04",
   492 => x"02fc050d",
   493 => x"8fba048c",
   494 => x"872d80f6",
   495 => x"518dbe2d",
   496 => x"bbdc08f3",
   497 => x"3880da51",
   498 => x"8dbe2dbb",
   499 => x"dc08e838",
   500 => x"bbdc08ba",
   501 => x"9c0cbbdc",
   502 => x"085184f0",
   503 => x"2d028405",
   504 => x"0d0402ec",
   505 => x"050d7654",
   506 => x"8052870b",
   507 => x"881580f5",
   508 => x"2d565374",
   509 => x"72248338",
   510 => x"a0537251",
   511 => x"82f92d81",
   512 => x"128b1580",
   513 => x"f52d5452",
   514 => x"727225de",
   515 => x"38029405",
   516 => x"0d0402f0",
   517 => x"050dbcb0",
   518 => x"085481f8",
   519 => x"2d800bbc",
   520 => x"b40c7308",
   521 => x"802e8180",
   522 => x"38820bbb",
   523 => x"f00cbcb4",
   524 => x"088f06bb",
   525 => x"ec0c7308",
   526 => x"5271832e",
   527 => x"96387183",
   528 => x"26893871",
   529 => x"812eaf38",
   530 => x"91930471",
   531 => x"852e9f38",
   532 => x"91930488",
   533 => x"1480f52d",
   534 => x"841508b5",
   535 => x"f0535452",
   536 => x"85fe2d71",
   537 => x"84291370",
   538 => x"08525291",
   539 => x"97047351",
   540 => x"8fe22d91",
   541 => x"9304ba98",
   542 => x"08881508",
   543 => x"2c708106",
   544 => x"51527180",
   545 => x"2e8738b5",
   546 => x"f4519190",
   547 => x"04b5f851",
   548 => x"85fe2d84",
   549 => x"14085185",
   550 => x"fe2dbcb4",
   551 => x"088105bc",
   552 => x"b40c8c14",
   553 => x"5490a204",
   554 => x"0290050d",
   555 => x"0471bcb0",
   556 => x"0c90922d",
   557 => x"bcb408ff",
   558 => x"05bcb80c",
   559 => x"0402e805",
   560 => x"0dbcb008",
   561 => x"bcbc0857",
   562 => x"5587518d",
   563 => x"be2dbbdc",
   564 => x"08812a70",
   565 => x"81065152",
   566 => x"71802ea0",
   567 => x"3891e304",
   568 => x"8c872d87",
   569 => x"518dbe2d",
   570 => x"bbdc08f4",
   571 => x"38ba9c08",
   572 => x"813270ba",
   573 => x"9c0c7052",
   574 => x"5284f02d",
   575 => x"80fe518d",
   576 => x"be2dbbdc",
   577 => x"08802ea6",
   578 => x"38ba9c08",
   579 => x"802e9138",
   580 => x"800bba9c",
   581 => x"0c805184",
   582 => x"f02d92a0",
   583 => x"048c872d",
   584 => x"80fe518d",
   585 => x"be2dbbdc",
   586 => x"08f33886",
   587 => x"f72dba9c",
   588 => x"08903881",
   589 => x"fd518dbe",
   590 => x"2d81fa51",
   591 => x"8dbe2d97",
   592 => x"f30481f5",
   593 => x"518dbe2d",
   594 => x"bbdc0881",
   595 => x"2a708106",
   596 => x"51527180",
   597 => x"2eaf38bc",
   598 => x"b8085271",
   599 => x"802e8938",
   600 => x"ff12bcb8",
   601 => x"0c938504",
   602 => x"bcb40810",
   603 => x"bcb40805",
   604 => x"70842916",
   605 => x"51528812",
   606 => x"08802e89",
   607 => x"38ff5188",
   608 => x"12085271",
   609 => x"2d81f251",
   610 => x"8dbe2dbb",
   611 => x"dc08812a",
   612 => x"70810651",
   613 => x"5271802e",
   614 => x"b138bcb4",
   615 => x"08ff11bc",
   616 => x"b8085653",
   617 => x"53737225",
   618 => x"89388114",
   619 => x"bcb80c93",
   620 => x"ca047210",
   621 => x"13708429",
   622 => x"16515288",
   623 => x"1208802e",
   624 => x"8938fe51",
   625 => x"88120852",
   626 => x"712d81fd",
   627 => x"518dbe2d",
   628 => x"bbdc0881",
   629 => x"2a708106",
   630 => x"51527180",
   631 => x"2ead38bc",
   632 => x"b808802e",
   633 => x"8938800b",
   634 => x"bcb80c94",
   635 => x"8b04bcb4",
   636 => x"0810bcb4",
   637 => x"08057084",
   638 => x"29165152",
   639 => x"88120880",
   640 => x"2e8938fd",
   641 => x"51881208",
   642 => x"52712d81",
   643 => x"fa518dbe",
   644 => x"2dbbdc08",
   645 => x"812a7081",
   646 => x"06515271",
   647 => x"802eae38",
   648 => x"bcb408ff",
   649 => x"115452bc",
   650 => x"b8087325",
   651 => x"883872bc",
   652 => x"b80c94cd",
   653 => x"04711012",
   654 => x"70842916",
   655 => x"51528812",
   656 => x"08802e89",
   657 => x"38fc5188",
   658 => x"12085271",
   659 => x"2dbcb808",
   660 => x"70535473",
   661 => x"802e8a38",
   662 => x"8c15ff15",
   663 => x"555594d3",
   664 => x"04820bbb",
   665 => x"f00c718f",
   666 => x"06bbec0c",
   667 => x"81eb518d",
   668 => x"be2dbbdc",
   669 => x"08812a70",
   670 => x"81065152",
   671 => x"71802ead",
   672 => x"38740885",
   673 => x"2e098106",
   674 => x"a4388815",
   675 => x"80f52dff",
   676 => x"05527188",
   677 => x"1681b72d",
   678 => x"71982b52",
   679 => x"71802588",
   680 => x"38800b88",
   681 => x"1681b72d",
   682 => x"74518fe2",
   683 => x"2d81f451",
   684 => x"8dbe2dbb",
   685 => x"dc08812a",
   686 => x"70810651",
   687 => x"5271802e",
   688 => x"b3387408",
   689 => x"852e0981",
   690 => x"06aa3888",
   691 => x"1580f52d",
   692 => x"81055271",
   693 => x"881681b7",
   694 => x"2d7181ff",
   695 => x"068b1680",
   696 => x"f52d5452",
   697 => x"72722787",
   698 => x"38728816",
   699 => x"81b72d74",
   700 => x"518fe22d",
   701 => x"80da518d",
   702 => x"be2dbbdc",
   703 => x"08812a70",
   704 => x"81065152",
   705 => x"71802e81",
   706 => x"a638bcb0",
   707 => x"08bcb808",
   708 => x"55537380",
   709 => x"2e8a388c",
   710 => x"13ff1555",
   711 => x"53969204",
   712 => x"72085271",
   713 => x"822ea638",
   714 => x"71822689",
   715 => x"3871812e",
   716 => x"a93897af",
   717 => x"0471832e",
   718 => x"b1387184",
   719 => x"2e098106",
   720 => x"80ed3888",
   721 => x"13085191",
   722 => x"ad2d97af",
   723 => x"04bcb808",
   724 => x"51881308",
   725 => x"52712d97",
   726 => x"af04810b",
   727 => x"8814082b",
   728 => x"ba980832",
   729 => x"ba980c97",
   730 => x"85048813",
   731 => x"80f52d81",
   732 => x"058b1480",
   733 => x"f52d5354",
   734 => x"71742483",
   735 => x"38805473",
   736 => x"881481b7",
   737 => x"2d90922d",
   738 => x"97af0475",
   739 => x"08802ea2",
   740 => x"38750851",
   741 => x"8dbe2dbb",
   742 => x"dc088106",
   743 => x"5271802e",
   744 => x"8b38bcb8",
   745 => x"08518416",
   746 => x"0852712d",
   747 => x"88165675",
   748 => x"da388054",
   749 => x"800bbbf0",
   750 => x"0c738f06",
   751 => x"bbec0ca0",
   752 => x"5273bcb8",
   753 => x"082e0981",
   754 => x"069838bc",
   755 => x"b408ff05",
   756 => x"74327009",
   757 => x"81057072",
   758 => x"079f2a91",
   759 => x"71315151",
   760 => x"53537151",
   761 => x"82f92d81",
   762 => x"14548e74",
   763 => x"25c638ba",
   764 => x"9c085271",
   765 => x"bbdc0c02",
   766 => x"98050d04",
   767 => x"02f4050d",
   768 => x"d45281ff",
   769 => x"720c7108",
   770 => x"5381ff72",
   771 => x"0c72882b",
   772 => x"83fe8006",
   773 => x"72087081",
   774 => x"ff065152",
   775 => x"5381ff72",
   776 => x"0c727107",
   777 => x"882b7208",
   778 => x"7081ff06",
   779 => x"51525381",
   780 => x"ff720c72",
   781 => x"7107882b",
   782 => x"72087081",
   783 => x"ff067207",
   784 => x"bbdc0c52",
   785 => x"53028c05",
   786 => x"0d0402f4",
   787 => x"050d7476",
   788 => x"7181ff06",
   789 => x"d40c5353",
   790 => x"bcc00885",
   791 => x"3871892b",
   792 => x"5271982a",
   793 => x"d40c7190",
   794 => x"2a7081ff",
   795 => x"06d40c51",
   796 => x"71882a70",
   797 => x"81ff06d4",
   798 => x"0c517181",
   799 => x"ff06d40c",
   800 => x"72902a70",
   801 => x"81ff06d4",
   802 => x"0c51d408",
   803 => x"7081ff06",
   804 => x"515182b8",
   805 => x"bf527081",
   806 => x"ff2e0981",
   807 => x"06943881",
   808 => x"ff0bd40c",
   809 => x"d4087081",
   810 => x"ff06ff14",
   811 => x"54515171",
   812 => x"e53870bb",
   813 => x"dc0c028c",
   814 => x"050d0402",
   815 => x"fc050d81",
   816 => x"c75181ff",
   817 => x"0bd40cff",
   818 => x"11517080",
   819 => x"25f43802",
   820 => x"84050d04",
   821 => x"02f4050d",
   822 => x"81ff0bd4",
   823 => x"0c935380",
   824 => x"5287fc80",
   825 => x"c15198ca",
   826 => x"2dbbdc08",
   827 => x"8b3881ff",
   828 => x"0bd40c81",
   829 => x"539a8104",
   830 => x"99bb2dff",
   831 => x"135372df",
   832 => x"3872bbdc",
   833 => x"0c028c05",
   834 => x"0d0402ec",
   835 => x"050d810b",
   836 => x"bcc00c84",
   837 => x"54d00870",
   838 => x"8f2a7081",
   839 => x"06515153",
   840 => x"72f33872",
   841 => x"d00c99bb",
   842 => x"2db5fc51",
   843 => x"85fe2dd0",
   844 => x"08708f2a",
   845 => x"70810651",
   846 => x"515372f3",
   847 => x"38810bd0",
   848 => x"0cb15380",
   849 => x"5284d480",
   850 => x"c05198ca",
   851 => x"2dbbdc08",
   852 => x"812e9338",
   853 => x"72822ebd",
   854 => x"38ff1353",
   855 => x"72e538ff",
   856 => x"145473ff",
   857 => x"b03899bb",
   858 => x"2d83aa52",
   859 => x"849c80c8",
   860 => x"5198ca2d",
   861 => x"bbdc0881",
   862 => x"2e098106",
   863 => x"923897fc",
   864 => x"2dbbdc08",
   865 => x"83ffff06",
   866 => x"537283aa",
   867 => x"2e9d3899",
   868 => x"d42d9ba6",
   869 => x"04b68851",
   870 => x"85fe2d80",
   871 => x"539cf404",
   872 => x"b6a05185",
   873 => x"fe2d8054",
   874 => x"9cc60481",
   875 => x"ff0bd40c",
   876 => x"b15499bb",
   877 => x"2d8fcf53",
   878 => x"805287fc",
   879 => x"80f75198",
   880 => x"ca2dbbdc",
   881 => x"0855bbdc",
   882 => x"08812e09",
   883 => x"81069b38",
   884 => x"81ff0bd4",
   885 => x"0c820a52",
   886 => x"849c80e9",
   887 => x"5198ca2d",
   888 => x"bbdc0880",
   889 => x"2e8d3899",
   890 => x"bb2dff13",
   891 => x"5372c938",
   892 => x"9cb90481",
   893 => x"ff0bd40c",
   894 => x"bbdc0852",
   895 => x"87fc80fa",
   896 => x"5198ca2d",
   897 => x"bbdc08b1",
   898 => x"3881ff0b",
   899 => x"d40cd408",
   900 => x"5381ff0b",
   901 => x"d40c81ff",
   902 => x"0bd40c81",
   903 => x"ff0bd40c",
   904 => x"81ff0bd4",
   905 => x"0c72862a",
   906 => x"70810676",
   907 => x"56515372",
   908 => x"9538bbdc",
   909 => x"08549cc6",
   910 => x"0473822e",
   911 => x"fee238ff",
   912 => x"145473fe",
   913 => x"ed3873bc",
   914 => x"c00c738b",
   915 => x"38815287",
   916 => x"fc80d051",
   917 => x"98ca2d81",
   918 => x"ff0bd40c",
   919 => x"d008708f",
   920 => x"2a708106",
   921 => x"51515372",
   922 => x"f33872d0",
   923 => x"0c81ff0b",
   924 => x"d40c8153",
   925 => x"72bbdc0c",
   926 => x"0294050d",
   927 => x"0402e805",
   928 => x"0d785580",
   929 => x"5681ff0b",
   930 => x"d40cd008",
   931 => x"708f2a70",
   932 => x"81065151",
   933 => x"5372f338",
   934 => x"82810bd0",
   935 => x"0c81ff0b",
   936 => x"d40c7752",
   937 => x"87fc80d1",
   938 => x"5198ca2d",
   939 => x"80dbc6df",
   940 => x"54bbdc08",
   941 => x"802e8a38",
   942 => x"b6c05185",
   943 => x"fe2d9e94",
   944 => x"0481ff0b",
   945 => x"d40cd408",
   946 => x"7081ff06",
   947 => x"51537281",
   948 => x"fe2e0981",
   949 => x"069d3880",
   950 => x"ff5397fc",
   951 => x"2dbbdc08",
   952 => x"75708405",
   953 => x"570cff13",
   954 => x"53728025",
   955 => x"ed388156",
   956 => x"9df904ff",
   957 => x"145473c9",
   958 => x"3881ff0b",
   959 => x"d40c81ff",
   960 => x"0bd40cd0",
   961 => x"08708f2a",
   962 => x"70810651",
   963 => x"515372f3",
   964 => x"3872d00c",
   965 => x"75bbdc0c",
   966 => x"0298050d",
   967 => x"0402e805",
   968 => x"0d77797b",
   969 => x"58555580",
   970 => x"53727625",
   971 => x"a3387470",
   972 => x"81055680",
   973 => x"f52d7470",
   974 => x"81055680",
   975 => x"f52d5252",
   976 => x"71712e86",
   977 => x"3881519e",
   978 => x"d2048113",
   979 => x"539ea904",
   980 => x"805170bb",
   981 => x"dc0c0298",
   982 => x"050d0402",
   983 => x"ec050d76",
   984 => x"5574802e",
   985 => x"be389a15",
   986 => x"80e02d51",
   987 => x"ac9f2dbb",
   988 => x"dc08bbdc",
   989 => x"0880c2f4",
   990 => x"0cbbdc08",
   991 => x"545480c2",
   992 => x"d008802e",
   993 => x"99389415",
   994 => x"80e02d51",
   995 => x"ac9f2dbb",
   996 => x"dc08902b",
   997 => x"83fff00a",
   998 => x"06707507",
   999 => x"51537280",
  1000 => x"c2f40c80",
  1001 => x"c2f40853",
  1002 => x"72802e9d",
  1003 => x"3880c2c8",
  1004 => x"08fe1471",
  1005 => x"2980c2dc",
  1006 => x"080580c2",
  1007 => x"f80c7084",
  1008 => x"2b80c2d4",
  1009 => x"0c549ff7",
  1010 => x"0480c2e0",
  1011 => x"0880c2f4",
  1012 => x"0c80c2e4",
  1013 => x"0880c2f8",
  1014 => x"0c80c2d0",
  1015 => x"08802e8b",
  1016 => x"3880c2c8",
  1017 => x"08842b53",
  1018 => x"9ff20480",
  1019 => x"c2e80884",
  1020 => x"2b537280",
  1021 => x"c2d40c02",
  1022 => x"94050d04",
  1023 => x"02d8050d",
  1024 => x"800b80c2",
  1025 => x"d00c8454",
  1026 => x"9a8a2dbb",
  1027 => x"dc08802e",
  1028 => x"9538bcc4",
  1029 => x"5280519c",
  1030 => x"fd2dbbdc",
  1031 => x"08802e86",
  1032 => x"38fe54a0",
  1033 => x"ae04ff14",
  1034 => x"54738024",
  1035 => x"db38738c",
  1036 => x"38b6d051",
  1037 => x"85fe2d73",
  1038 => x"55a5d804",
  1039 => x"8056810b",
  1040 => x"80c2fc0c",
  1041 => x"8853b6e4",
  1042 => x"52bcfa51",
  1043 => x"9e9d2dbb",
  1044 => x"dc08762e",
  1045 => x"09810688",
  1046 => x"38bbdc08",
  1047 => x"80c2fc0c",
  1048 => x"8853b6f0",
  1049 => x"52bd9651",
  1050 => x"9e9d2dbb",
  1051 => x"dc088838",
  1052 => x"bbdc0880",
  1053 => x"c2fc0c80",
  1054 => x"c2fc0880",
  1055 => x"2e80fc38",
  1056 => x"80c08a0b",
  1057 => x"80f52d80",
  1058 => x"c08b0b80",
  1059 => x"f52d7198",
  1060 => x"2b71902b",
  1061 => x"0780c08c",
  1062 => x"0b80f52d",
  1063 => x"70882b72",
  1064 => x"0780c08d",
  1065 => x"0b80f52d",
  1066 => x"710780c0",
  1067 => x"c20b80f5",
  1068 => x"2d80c0c3",
  1069 => x"0b80f52d",
  1070 => x"71882b07",
  1071 => x"535f5452",
  1072 => x"5a565755",
  1073 => x"7381abaa",
  1074 => x"2e098106",
  1075 => x"8d387551",
  1076 => x"abef2dbb",
  1077 => x"dc0856a1",
  1078 => x"e7047382",
  1079 => x"d4d52e87",
  1080 => x"38b6fc51",
  1081 => x"a2a904bc",
  1082 => x"c4527551",
  1083 => x"9cfd2dbb",
  1084 => x"dc0855bb",
  1085 => x"dc08802e",
  1086 => x"83de3888",
  1087 => x"53b6f052",
  1088 => x"bd96519e",
  1089 => x"9d2dbbdc",
  1090 => x"088a3881",
  1091 => x"0b80c2d0",
  1092 => x"0ca2af04",
  1093 => x"8853b6e4",
  1094 => x"52bcfa51",
  1095 => x"9e9d2dbb",
  1096 => x"dc08802e",
  1097 => x"8a38b790",
  1098 => x"5185fe2d",
  1099 => x"a38b0480",
  1100 => x"c0c20b80",
  1101 => x"f52d5473",
  1102 => x"80d52e09",
  1103 => x"810680cb",
  1104 => x"3880c0c3",
  1105 => x"0b80f52d",
  1106 => x"547381aa",
  1107 => x"2e098106",
  1108 => x"ba38800b",
  1109 => x"bcc40b80",
  1110 => x"f52d5654",
  1111 => x"7481e92e",
  1112 => x"83388154",
  1113 => x"7481eb2e",
  1114 => x"8c388055",
  1115 => x"73752e09",
  1116 => x"810682e4",
  1117 => x"38bccf0b",
  1118 => x"80f52d55",
  1119 => x"748d38bc",
  1120 => x"d00b80f5",
  1121 => x"2d547382",
  1122 => x"2e863880",
  1123 => x"55a5d804",
  1124 => x"bcd10b80",
  1125 => x"f52d7080",
  1126 => x"c2c80cff",
  1127 => x"0580c2cc",
  1128 => x"0cbcd20b",
  1129 => x"80f52dbc",
  1130 => x"d30b80f5",
  1131 => x"2d587605",
  1132 => x"77828029",
  1133 => x"057080c2",
  1134 => x"d80cbcd4",
  1135 => x"0b80f52d",
  1136 => x"7080c2ec",
  1137 => x"0c80c2d0",
  1138 => x"08595758",
  1139 => x"76802e81",
  1140 => x"ac388853",
  1141 => x"b6f052bd",
  1142 => x"96519e9d",
  1143 => x"2dbbdc08",
  1144 => x"81f63880",
  1145 => x"c2c80870",
  1146 => x"842b80c2",
  1147 => x"d40c7080",
  1148 => x"c2e80cbc",
  1149 => x"e90b80f5",
  1150 => x"2dbce80b",
  1151 => x"80f52d71",
  1152 => x"82802905",
  1153 => x"bcea0b80",
  1154 => x"f52d7084",
  1155 => x"80802912",
  1156 => x"bceb0b80",
  1157 => x"f52d7081",
  1158 => x"800a2912",
  1159 => x"7080c2f0",
  1160 => x"0c80c2ec",
  1161 => x"08712980",
  1162 => x"c2d80805",
  1163 => x"7080c2dc",
  1164 => x"0cbcf10b",
  1165 => x"80f52dbc",
  1166 => x"f00b80f5",
  1167 => x"2d718280",
  1168 => x"2905bcf2",
  1169 => x"0b80f52d",
  1170 => x"70848080",
  1171 => x"2912bcf3",
  1172 => x"0b80f52d",
  1173 => x"70982b81",
  1174 => x"f00a0672",
  1175 => x"057080c2",
  1176 => x"e00cfe11",
  1177 => x"7e297705",
  1178 => x"80c2e40c",
  1179 => x"52595243",
  1180 => x"545e5152",
  1181 => x"59525d57",
  1182 => x"5957a5d1",
  1183 => x"04bcd60b",
  1184 => x"80f52dbc",
  1185 => x"d50b80f5",
  1186 => x"2d718280",
  1187 => x"29057080",
  1188 => x"c2d40c70",
  1189 => x"a02983ff",
  1190 => x"0570892a",
  1191 => x"7080c2e8",
  1192 => x"0cbcdb0b",
  1193 => x"80f52dbc",
  1194 => x"da0b80f5",
  1195 => x"2d718280",
  1196 => x"29057080",
  1197 => x"c2f00c7b",
  1198 => x"71291e70",
  1199 => x"80c2e40c",
  1200 => x"7d80c2e0",
  1201 => x"0c730580",
  1202 => x"c2dc0c55",
  1203 => x"5e515155",
  1204 => x"5580519e",
  1205 => x"db2d8155",
  1206 => x"74bbdc0c",
  1207 => x"02a8050d",
  1208 => x"0402ec05",
  1209 => x"0d767087",
  1210 => x"2c7180ff",
  1211 => x"06555654",
  1212 => x"80c2d008",
  1213 => x"8a387388",
  1214 => x"2c7481ff",
  1215 => x"065455bc",
  1216 => x"c45280c2",
  1217 => x"d8081551",
  1218 => x"9cfd2dbb",
  1219 => x"dc0854bb",
  1220 => x"dc08802e",
  1221 => x"b43880c2",
  1222 => x"d008802e",
  1223 => x"98387284",
  1224 => x"29bcc405",
  1225 => x"70085253",
  1226 => x"abef2dbb",
  1227 => x"dc08f00a",
  1228 => x"0653a6c7",
  1229 => x"047210bc",
  1230 => x"c4057080",
  1231 => x"e02d5253",
  1232 => x"ac9f2dbb",
  1233 => x"dc085372",
  1234 => x"5473bbdc",
  1235 => x"0c029405",
  1236 => x"0d0402e0",
  1237 => x"050d7970",
  1238 => x"842c80c2",
  1239 => x"f8080571",
  1240 => x"8f065255",
  1241 => x"53728938",
  1242 => x"bcc45273",
  1243 => x"519cfd2d",
  1244 => x"72a029bc",
  1245 => x"c4055480",
  1246 => x"7480f52d",
  1247 => x"56537473",
  1248 => x"2e833881",
  1249 => x"537481e5",
  1250 => x"2e81f138",
  1251 => x"81707406",
  1252 => x"54587280",
  1253 => x"2e81e538",
  1254 => x"8b1480f5",
  1255 => x"2d70832a",
  1256 => x"79065856",
  1257 => x"769938ba",
  1258 => x"a0085372",
  1259 => x"89387280",
  1260 => x"c0c40b81",
  1261 => x"b72d76ba",
  1262 => x"a00c7353",
  1263 => x"a8fe0475",
  1264 => x"8f2e0981",
  1265 => x"0681b538",
  1266 => x"749f068d",
  1267 => x"2980c0b7",
  1268 => x"11515381",
  1269 => x"1480f52d",
  1270 => x"73708105",
  1271 => x"5581b72d",
  1272 => x"831480f5",
  1273 => x"2d737081",
  1274 => x"055581b7",
  1275 => x"2d851480",
  1276 => x"f52d7370",
  1277 => x"81055581",
  1278 => x"b72d8714",
  1279 => x"80f52d73",
  1280 => x"70810555",
  1281 => x"81b72d89",
  1282 => x"1480f52d",
  1283 => x"73708105",
  1284 => x"5581b72d",
  1285 => x"8e1480f5",
  1286 => x"2d737081",
  1287 => x"055581b7",
  1288 => x"2d901480",
  1289 => x"f52d7370",
  1290 => x"81055581",
  1291 => x"b72d9214",
  1292 => x"80f52d73",
  1293 => x"70810555",
  1294 => x"81b72d94",
  1295 => x"1480f52d",
  1296 => x"73708105",
  1297 => x"5581b72d",
  1298 => x"961480f5",
  1299 => x"2d737081",
  1300 => x"055581b7",
  1301 => x"2d981480",
  1302 => x"f52d7370",
  1303 => x"81055581",
  1304 => x"b72d9c14",
  1305 => x"80f52d73",
  1306 => x"70810555",
  1307 => x"81b72d9e",
  1308 => x"1480f52d",
  1309 => x"7381b72d",
  1310 => x"77baa00c",
  1311 => x"805372bb",
  1312 => x"dc0c02a0",
  1313 => x"050d0402",
  1314 => x"cc050d7e",
  1315 => x"605e5a80",
  1316 => x"0b80c2f4",
  1317 => x"0880c2f8",
  1318 => x"08595c56",
  1319 => x"805880c2",
  1320 => x"d408782e",
  1321 => x"81b03877",
  1322 => x"8f06a017",
  1323 => x"5754738f",
  1324 => x"38bcc452",
  1325 => x"76518117",
  1326 => x"579cfd2d",
  1327 => x"bcc45680",
  1328 => x"7680f52d",
  1329 => x"56547474",
  1330 => x"2e833881",
  1331 => x"547481e5",
  1332 => x"2e80f738",
  1333 => x"81707506",
  1334 => x"555c7380",
  1335 => x"2e80eb38",
  1336 => x"8b1680f5",
  1337 => x"2d980659",
  1338 => x"7880df38",
  1339 => x"8b537c52",
  1340 => x"75519e9d",
  1341 => x"2dbbdc08",
  1342 => x"80d0389c",
  1343 => x"160851ab",
  1344 => x"ef2dbbdc",
  1345 => x"08841b0c",
  1346 => x"9a1680e0",
  1347 => x"2d51ac9f",
  1348 => x"2dbbdc08",
  1349 => x"bbdc0888",
  1350 => x"1c0cbbdc",
  1351 => x"08555580",
  1352 => x"c2d00880",
  1353 => x"2e983894",
  1354 => x"1680e02d",
  1355 => x"51ac9f2d",
  1356 => x"bbdc0890",
  1357 => x"2b83fff0",
  1358 => x"0a067016",
  1359 => x"51547388",
  1360 => x"1b0c787a",
  1361 => x"0c7b54ab",
  1362 => x"8f048118",
  1363 => x"5880c2d4",
  1364 => x"087826fe",
  1365 => x"d23880c2",
  1366 => x"d008802e",
  1367 => x"b0387a51",
  1368 => x"a5e12dbb",
  1369 => x"dc08bbdc",
  1370 => x"0880ffff",
  1371 => x"fff80655",
  1372 => x"5b7380ff",
  1373 => x"fffff82e",
  1374 => x"9438bbdc",
  1375 => x"08fe0580",
  1376 => x"c2c80829",
  1377 => x"80c2dc08",
  1378 => x"0557a99c",
  1379 => x"04805473",
  1380 => x"bbdc0c02",
  1381 => x"b4050d04",
  1382 => x"02f4050d",
  1383 => x"74700881",
  1384 => x"05710c70",
  1385 => x"0880c2cc",
  1386 => x"08065353",
  1387 => x"718e3888",
  1388 => x"130851a5",
  1389 => x"e12dbbdc",
  1390 => x"0888140c",
  1391 => x"810bbbdc",
  1392 => x"0c028c05",
  1393 => x"0d0402f0",
  1394 => x"050d7588",
  1395 => x"1108fe05",
  1396 => x"80c2c808",
  1397 => x"2980c2dc",
  1398 => x"08117208",
  1399 => x"80c2cc08",
  1400 => x"06057955",
  1401 => x"5354549c",
  1402 => x"fd2d0290",
  1403 => x"050d0402",
  1404 => x"f4050d74",
  1405 => x"70882a83",
  1406 => x"fe800670",
  1407 => x"72982a07",
  1408 => x"72882b87",
  1409 => x"fc808006",
  1410 => x"73982b81",
  1411 => x"f00a0671",
  1412 => x"730707bb",
  1413 => x"dc0c5651",
  1414 => x"5351028c",
  1415 => x"050d0402",
  1416 => x"f8050d02",
  1417 => x"8e0580f5",
  1418 => x"2d74882b",
  1419 => x"077083ff",
  1420 => x"ff06bbdc",
  1421 => x"0c510288",
  1422 => x"050d0402",
  1423 => x"f4050d74",
  1424 => x"76785354",
  1425 => x"52807125",
  1426 => x"97387270",
  1427 => x"81055480",
  1428 => x"f52d7270",
  1429 => x"81055481",
  1430 => x"b72dff11",
  1431 => x"5170eb38",
  1432 => x"807281b7",
  1433 => x"2d028c05",
  1434 => x"0d0402e8",
  1435 => x"050d7756",
  1436 => x"80705654",
  1437 => x"737624b3",
  1438 => x"3880c2d4",
  1439 => x"08742eab",
  1440 => x"387351a6",
  1441 => x"d22dbbdc",
  1442 => x"08bbdc08",
  1443 => x"09810570",
  1444 => x"bbdc0807",
  1445 => x"9f2a7705",
  1446 => x"81175757",
  1447 => x"53537476",
  1448 => x"24893880",
  1449 => x"c2d40874",
  1450 => x"26d73872",
  1451 => x"bbdc0c02",
  1452 => x"98050d04",
  1453 => x"02f0050d",
  1454 => x"bbd80816",
  1455 => x"51acea2d",
  1456 => x"bbdc0880",
  1457 => x"2e9e388b",
  1458 => x"53bbdc08",
  1459 => x"5280c0c4",
  1460 => x"51acbb2d",
  1461 => x"80c38008",
  1462 => x"5473802e",
  1463 => x"873880c0",
  1464 => x"c451732d",
  1465 => x"0290050d",
  1466 => x"0402dc05",
  1467 => x"0d80705a",
  1468 => x"5574bbd8",
  1469 => x"0825b138",
  1470 => x"80c2d408",
  1471 => x"752ea938",
  1472 => x"7851a6d2",
  1473 => x"2dbbdc08",
  1474 => x"09810570",
  1475 => x"bbdc0807",
  1476 => x"9f2a7605",
  1477 => x"811b5b56",
  1478 => x"5474bbd8",
  1479 => x"08258938",
  1480 => x"80c2d408",
  1481 => x"7926d938",
  1482 => x"80557880",
  1483 => x"c2d40827",
  1484 => x"81d43878",
  1485 => x"51a6d22d",
  1486 => x"bbdc0880",
  1487 => x"2e81a838",
  1488 => x"bbdc088b",
  1489 => x"0580f52d",
  1490 => x"70842a70",
  1491 => x"81067710",
  1492 => x"78842b80",
  1493 => x"c0c40b80",
  1494 => x"f52d5c5c",
  1495 => x"53515556",
  1496 => x"73802e80",
  1497 => x"c9387416",
  1498 => x"822bb0aa",
  1499 => x"0bbaac12",
  1500 => x"0c547775",
  1501 => x"311080c3",
  1502 => x"84115556",
  1503 => x"90747081",
  1504 => x"055681b7",
  1505 => x"2da07481",
  1506 => x"b72d7681",
  1507 => x"ff068116",
  1508 => x"58547380",
  1509 => x"2e8a389c",
  1510 => x"5380c0c4",
  1511 => x"52afa604",
  1512 => x"8b53bbdc",
  1513 => x"085280c3",
  1514 => x"861651af",
  1515 => x"df047416",
  1516 => x"822badb4",
  1517 => x"0bbaac12",
  1518 => x"0c547681",
  1519 => x"ff068116",
  1520 => x"58547380",
  1521 => x"2e8a389c",
  1522 => x"5380c0c4",
  1523 => x"52afd604",
  1524 => x"8b53bbdc",
  1525 => x"08527775",
  1526 => x"311080c3",
  1527 => x"84055176",
  1528 => x"55acbb2d",
  1529 => x"affb0474",
  1530 => x"90297531",
  1531 => x"701080c3",
  1532 => x"84055154",
  1533 => x"bbdc0874",
  1534 => x"81b72d81",
  1535 => x"1959748b",
  1536 => x"24a338ae",
  1537 => x"aa047490",
  1538 => x"29753170",
  1539 => x"1080c384",
  1540 => x"058c7731",
  1541 => x"57515480",
  1542 => x"7481b72d",
  1543 => x"9e14ff16",
  1544 => x"565474f3",
  1545 => x"3802a405",
  1546 => x"0d0402fc",
  1547 => x"050dbbd8",
  1548 => x"081351ac",
  1549 => x"ea2dbbdc",
  1550 => x"08802e88",
  1551 => x"38bbdc08",
  1552 => x"519edb2d",
  1553 => x"800bbbd8",
  1554 => x"0cade92d",
  1555 => x"90922d02",
  1556 => x"84050d04",
  1557 => x"02fc050d",
  1558 => x"725170fd",
  1559 => x"2ead3870",
  1560 => x"fd248a38",
  1561 => x"70fc2e80",
  1562 => x"c438b1b5",
  1563 => x"0470fe2e",
  1564 => x"b13870ff",
  1565 => x"2e098106",
  1566 => x"bc38bbd8",
  1567 => x"08517080",
  1568 => x"2eb338ff",
  1569 => x"11bbd80c",
  1570 => x"b1b504bb",
  1571 => x"d808f005",
  1572 => x"70bbd80c",
  1573 => x"51708025",
  1574 => x"9c38800b",
  1575 => x"bbd80cb1",
  1576 => x"b504bbd8",
  1577 => x"088105bb",
  1578 => x"d80cb1b5",
  1579 => x"04bbd808",
  1580 => x"9005bbd8",
  1581 => x"0cade92d",
  1582 => x"90922d02",
  1583 => x"84050d04",
  1584 => x"02fc050d",
  1585 => x"800bbbd8",
  1586 => x"0cade92d",
  1587 => x"8fa92dbb",
  1588 => x"dc08bbc8",
  1589 => x"0cbaa451",
  1590 => x"91ad2d02",
  1591 => x"84050d04",
  1592 => x"7180c380",
  1593 => x"0c040000",
  1594 => x"00ffffff",
  1595 => x"ff00ffff",
  1596 => x"ffff00ff",
  1597 => x"ffffff00",
  1598 => x"52657365",
  1599 => x"74202620",
  1600 => x"536f6c74",
  1601 => x"61722043",
  1602 => x"61727475",
  1603 => x"63686f00",
  1604 => x"506c6179",
  1605 => x"2f53746f",
  1606 => x"70204369",
  1607 => x"6e746100",
  1608 => x"43617267",
  1609 => x"61722044",
  1610 => x"6973636f",
  1611 => x"2f43696e",
  1612 => x"74612f43",
  1613 => x"61727420",
  1614 => x"10000000",
  1615 => x"45786974",
  1616 => x"00000000",
  1617 => x"44697363",
  1618 => x"6f204772",
  1619 => x"61626162",
  1620 => x"6c650000",
  1621 => x"44697363",
  1622 => x"6f20536f",
  1623 => x"6c6f204c",
  1624 => x"65637475",
  1625 => x"72610000",
  1626 => x"50756572",
  1627 => x"746f2055",
  1628 => x"41525400",
  1629 => x"50756572",
  1630 => x"746f2034",
  1631 => x"20506c61",
  1632 => x"79657273",
  1633 => x"00000000",
  1634 => x"536f6e69",
  1635 => x"646f2043",
  1636 => x"696e7461",
  1637 => x"204f6666",
  1638 => x"00000000",
  1639 => x"536f6e69",
  1640 => x"646f2043",
  1641 => x"696e7461",
  1642 => x"204f6e00",
  1643 => x"4a6f7973",
  1644 => x"7469636b",
  1645 => x"73204e6f",
  1646 => x"726d616c",
  1647 => x"00000000",
  1648 => x"4a6f7973",
  1649 => x"7469636b",
  1650 => x"7320496e",
  1651 => x"74657263",
  1652 => x"616d6269",
  1653 => x"61646f73",
  1654 => x"00000000",
  1655 => x"41756469",
  1656 => x"6f204669",
  1657 => x"6c746572",
  1658 => x"204f6e00",
  1659 => x"41756469",
  1660 => x"6f204669",
  1661 => x"6c746572",
  1662 => x"204f6666",
  1663 => x"00000000",
  1664 => x"43494120",
  1665 => x"36323536",
  1666 => x"00000000",
  1667 => x"43494120",
  1668 => x"38353231",
  1669 => x"00000000",
  1670 => x"53494420",
  1671 => x"36353831",
  1672 => x"204d6f6e",
  1673 => x"6f000000",
  1674 => x"53494420",
  1675 => x"36353831",
  1676 => x"20537465",
  1677 => x"72656f00",
  1678 => x"53494420",
  1679 => x"38353830",
  1680 => x"204d6f6e",
  1681 => x"6f000000",
  1682 => x"53494420",
  1683 => x"38353830",
  1684 => x"20537465",
  1685 => x"72656f00",
  1686 => x"53494420",
  1687 => x"50736575",
  1688 => x"646f2053",
  1689 => x"74657265",
  1690 => x"6f000000",
  1691 => x"56696465",
  1692 => x"6f205041",
  1693 => x"4c000000",
  1694 => x"56696465",
  1695 => x"6f204e54",
  1696 => x"53430000",
  1697 => x"5363616e",
  1698 => x"6c696e65",
  1699 => x"73204e6f",
  1700 => x"6e650000",
  1701 => x"5363616e",
  1702 => x"6c696e65",
  1703 => x"73204352",
  1704 => x"54203235",
  1705 => x"25000000",
  1706 => x"5363616e",
  1707 => x"6c696e65",
  1708 => x"73204352",
  1709 => x"54203530",
  1710 => x"25000000",
  1711 => x"5363616e",
  1712 => x"6c696e65",
  1713 => x"73204352",
  1714 => x"54203735",
  1715 => x"25000000",
  1716 => x"43617267",
  1717 => x"61204661",
  1718 => x"6c6c6964",
  1719 => x"61000000",
  1720 => x"4f4b0000",
  1721 => x"43363420",
  1722 => x"20202020",
  1723 => x"44415400",
  1724 => x"16200000",
  1725 => x"14200000",
  1726 => x"15200000",
  1727 => x"53442069",
  1728 => x"6e69742e",
  1729 => x"2e2e0a00",
  1730 => x"53442063",
  1731 => x"61726420",
  1732 => x"72657365",
  1733 => x"74206661",
  1734 => x"696c6564",
  1735 => x"210a0000",
  1736 => x"53444843",
  1737 => x"20657272",
  1738 => x"6f72210a",
  1739 => x"00000000",
  1740 => x"57726974",
  1741 => x"65206661",
  1742 => x"696c6564",
  1743 => x"0a000000",
  1744 => x"52656164",
  1745 => x"20666169",
  1746 => x"6c65640a",
  1747 => x"00000000",
  1748 => x"43617264",
  1749 => x"20696e69",
  1750 => x"74206661",
  1751 => x"696c6564",
  1752 => x"0a000000",
  1753 => x"46415431",
  1754 => x"36202020",
  1755 => x"00000000",
  1756 => x"46415433",
  1757 => x"32202020",
  1758 => x"00000000",
  1759 => x"4e6f2070",
  1760 => x"61727469",
  1761 => x"74696f6e",
  1762 => x"20736967",
  1763 => x"0a000000",
  1764 => x"42616420",
  1765 => x"70617274",
  1766 => x"0a000000",
  1767 => x"4261636b",
  1768 => x"00000000",
  1769 => x"00000002",
  1770 => x"00000002",
  1771 => x"000018f8",
  1772 => x"0000034e",
  1773 => x"00000002",
  1774 => x"00001910",
  1775 => x"00000362",
  1776 => x"00000003",
  1777 => x"00001c9c",
  1778 => x"00000004",
  1779 => x"00000003",
  1780 => x"00001c94",
  1781 => x"00000002",
  1782 => x"00000003",
  1783 => x"00001c80",
  1784 => x"00000005",
  1785 => x"00000003",
  1786 => x"00001c78",
  1787 => x"00000002",
  1788 => x"00000003",
  1789 => x"00001c70",
  1790 => x"00000002",
  1791 => x"00000003",
  1792 => x"00001c68",
  1793 => x"00000002",
  1794 => x"00000003",
  1795 => x"00001c60",
  1796 => x"00000002",
  1797 => x"00000003",
  1798 => x"00001c58",
  1799 => x"00000002",
  1800 => x"00000003",
  1801 => x"00001c50",
  1802 => x"00000002",
  1803 => x"00000002",
  1804 => x"00001920",
  1805 => x"000018c0",
  1806 => x"00000002",
  1807 => x"0000193c",
  1808 => x"000007b0",
  1809 => x"00000000",
  1810 => x"00000000",
  1811 => x"00000000",
  1812 => x"00001944",
  1813 => x"00001954",
  1814 => x"00001968",
  1815 => x"00001974",
  1816 => x"00001988",
  1817 => x"0000199c",
  1818 => x"000019ac",
  1819 => x"000019c0",
  1820 => x"000019dc",
  1821 => x"000019ec",
  1822 => x"00001a00",
  1823 => x"00001a0c",
  1824 => x"00001a18",
  1825 => x"00001a28",
  1826 => x"00001a38",
  1827 => x"00001a48",
  1828 => x"00001a58",
  1829 => x"00001a6c",
  1830 => x"00001a78",
  1831 => x"00001a84",
  1832 => x"00001a94",
  1833 => x"00001aa8",
  1834 => x"00001abc",
  1835 => x"00000004",
  1836 => x"00001ad0",
  1837 => x"00001cac",
  1838 => x"00000004",
  1839 => x"00001ae0",
  1840 => x"00001ba8",
  1841 => x"00000000",
  1842 => x"00000000",
  1843 => x"00000000",
  1844 => x"00000000",
  1845 => x"00000000",
  1846 => x"00000000",
  1847 => x"00000000",
  1848 => x"00000000",
  1849 => x"00000000",
  1850 => x"00000000",
  1851 => x"00000000",
  1852 => x"00000000",
  1853 => x"00000000",
  1854 => x"00000000",
  1855 => x"00000000",
  1856 => x"00000000",
  1857 => x"00000000",
  1858 => x"00000000",
  1859 => x"00000000",
  1860 => x"00000000",
  1861 => x"00000000",
  1862 => x"00000000",
  1863 => x"00000000",
  1864 => x"00000000",
  1865 => x"00000002",
  1866 => x"00002184",
  1867 => x"000016b4",
  1868 => x"00000002",
  1869 => x"000021a2",
  1870 => x"000016b4",
  1871 => x"00000002",
  1872 => x"000021c0",
  1873 => x"000016b4",
  1874 => x"00000002",
  1875 => x"000021de",
  1876 => x"000016b4",
  1877 => x"00000002",
  1878 => x"000021fc",
  1879 => x"000016b4",
  1880 => x"00000002",
  1881 => x"0000221a",
  1882 => x"000016b4",
  1883 => x"00000002",
  1884 => x"00002238",
  1885 => x"000016b4",
  1886 => x"00000002",
  1887 => x"00002256",
  1888 => x"000016b4",
  1889 => x"00000002",
  1890 => x"00002274",
  1891 => x"000016b4",
  1892 => x"00000002",
  1893 => x"00002292",
  1894 => x"000016b4",
  1895 => x"00000002",
  1896 => x"000022b0",
  1897 => x"000016b4",
  1898 => x"00000002",
  1899 => x"000022ce",
  1900 => x"000016b4",
  1901 => x"00000002",
  1902 => x"000022ec",
  1903 => x"000016b4",
  1904 => x"00000004",
  1905 => x"00001b9c",
  1906 => x"00000000",
  1907 => x"00000000",
  1908 => x"00000000",
  1909 => x"00001854",
  1910 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

